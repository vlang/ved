module main

fn focus_app(next, event, data voidptr) {
	println('TODO: focus_app')
}

fn reg_key_vid() {
	println('TODO: reg_key_vid')
}


