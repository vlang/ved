module uiold

fn focus_app(next voidptr, event voidptr, data voidptr) {
}

pub fn reg_key_vid() {
}
