module uiold

fn focus_app(next voidptr, event voidptrs, data voidptr) {
}

pub fn reg_key_vid() {
}
